LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FOUR_BIT_COUNTER IS
	PORT(CLK : IN STD_LOGIC;
		  RST : IN STD_LOGIC;
		  BITS_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END FOUR_BIT_COUNTER;

ARCHITECTURE LOGIC OF FOUR_BIT_COUNTER IS
	SIGNAL COUNTER : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL WIRE : STD_LOGIC_vECTOR(5 DOWNTO 0) := (OTHERS => '0');
BEGIN
	WIRE(0) <= NOT COUNTER(3) AND COUNTER(2) AND COUNTER(1) AND COUNTER(0);
	WIRE(1) <= NOT COUNTER(2) OR NOT COUNTER(1) OR NOT COUNTER(0);
	WIRE(2) <= NOT COUNTER(1) OR NOT COUNTER(0);
	WIRE(3) <= NOT COUNTER(2) AND COUNTER(1) AND COUNTER(0);
	WIRE(4) <= COUNTER(3) AND WIRE(1);
	WIRE(5) <= COUNTER(2) AND WIRE(2);
	PROCESS(CLK, RST)
	BEGIN
		IF RST = '1' THEN
			COUNTER <= (OTHERS => '0');
		ELSIF CLK'EVENT AND CLK = '1' THEN
			COUNTER(3) <= WIRE(0) OR WIRE(4);
			COUNTER(2) <= WIRE(5) OR WIRE(3);
			COUNTER(1) <= COUNTER(1) XOR COUNTER(0);
			COUNTER(0) <= NOT COUNTER(0);
		END IF;
	END PROCESS;
	BITS_OUT(3 DOWNTO 0) <= COUNTER(3 DOWNTO 0);
END LOGIC;
		  